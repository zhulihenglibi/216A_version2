library verilog;
use verilog.vl_types.all;
entity adc_engine is
end adc_engine;
